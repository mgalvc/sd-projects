// processor.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module processor (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] nios_ii_data_master_readdata;                          // mm_interconnect_0:nios_II_data_master_readdata -> nios_II:d_readdata
	wire         nios_ii_data_master_waitrequest;                       // mm_interconnect_0:nios_II_data_master_waitrequest -> nios_II:d_waitrequest
	wire         nios_ii_data_master_debugaccess;                       // nios_II:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_II_data_master_debugaccess
	wire  [16:0] nios_ii_data_master_address;                           // nios_II:d_address -> mm_interconnect_0:nios_II_data_master_address
	wire   [3:0] nios_ii_data_master_byteenable;                        // nios_II:d_byteenable -> mm_interconnect_0:nios_II_data_master_byteenable
	wire         nios_ii_data_master_read;                              // nios_II:d_read -> mm_interconnect_0:nios_II_data_master_read
	wire         nios_ii_data_master_write;                             // nios_II:d_write -> mm_interconnect_0:nios_II_data_master_write
	wire  [31:0] nios_ii_data_master_writedata;                         // nios_II:d_writedata -> mm_interconnect_0:nios_II_data_master_writedata
	wire  [31:0] nios_ii_instruction_master_readdata;                   // mm_interconnect_0:nios_II_instruction_master_readdata -> nios_II:i_readdata
	wire         nios_ii_instruction_master_waitrequest;                // mm_interconnect_0:nios_II_instruction_master_waitrequest -> nios_II:i_waitrequest
	wire  [16:0] nios_ii_instruction_master_address;                    // nios_II:i_address -> mm_interconnect_0:nios_II_instruction_master_address
	wire         nios_ii_instruction_master_read;                       // nios_II:i_read -> mm_interconnect_0:nios_II_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios_ii_debug_mem_slave_readdata;    // nios_II:debug_mem_slave_readdata -> mm_interconnect_0:nios_II_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_waitrequest; // nios_II:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_II_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_debugaccess; // mm_interconnect_0:nios_II_debug_mem_slave_debugaccess -> nios_II:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_ii_debug_mem_slave_address;     // mm_interconnect_0:nios_II_debug_mem_slave_address -> nios_II:debug_mem_slave_address
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_read;        // mm_interconnect_0:nios_II_debug_mem_slave_read -> nios_II:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_ii_debug_mem_slave_byteenable;  // mm_interconnect_0:nios_II_debug_mem_slave_byteenable -> nios_II:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_write;       // mm_interconnect_0:nios_II_debug_mem_slave_write -> nios_II:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_ii_debug_mem_slave_writedata;   // mm_interconnect_0:nios_II_debug_mem_slave_writedata -> nios_II:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;                // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                  // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire  [12:0] mm_interconnect_0_memory_s1_address;                   // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                     // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                 // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                     // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire  [31:0] nios_ii_irq_irq;                                       // irq_mapper:sender_irq -> nios_II:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [irq_mapper:reset, memory:reset, mm_interconnect_0:nios_II_reset_reset_bridge_in_reset_reset, nios_II:reset_n]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [memory:reset_req, nios_II:reset_req, rst_translator:reset_req_in]
	wire         nios_ii_debug_reset_request_reset;                     // nios_II:debug_reset_request -> rst_controller:reset_in1

	custom_instruction custom_0 (
		.dataa  (), // nios_custom_instruction_slave.dataa
		.result ()  //                              .reset
	);

	processor_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	processor_nios_II nios_ii (
		.clk                                 (clk_clk),                                               //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (nios_ii_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_ii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_ii_data_master_read),                              //                          .read
		.d_readdata                          (nios_ii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_ii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_ii_data_master_write),                             //                          .write
		.d_writedata                         (nios_ii_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_ii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_ii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_ii_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_ii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_ii_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_ii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_ii_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_ii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_ii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_ii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_ii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_ii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_ii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_ii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_ii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	processor_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                               //                           clk_0_clk.clk
		.nios_II_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // nios_II_reset_reset_bridge_in_reset.reset
		.nios_II_data_master_address               (nios_ii_data_master_address),                           //                 nios_II_data_master.address
		.nios_II_data_master_waitrequest           (nios_ii_data_master_waitrequest),                       //                                    .waitrequest
		.nios_II_data_master_byteenable            (nios_ii_data_master_byteenable),                        //                                    .byteenable
		.nios_II_data_master_read                  (nios_ii_data_master_read),                              //                                    .read
		.nios_II_data_master_readdata              (nios_ii_data_master_readdata),                          //                                    .readdata
		.nios_II_data_master_write                 (nios_ii_data_master_write),                             //                                    .write
		.nios_II_data_master_writedata             (nios_ii_data_master_writedata),                         //                                    .writedata
		.nios_II_data_master_debugaccess           (nios_ii_data_master_debugaccess),                       //                                    .debugaccess
		.nios_II_instruction_master_address        (nios_ii_instruction_master_address),                    //          nios_II_instruction_master.address
		.nios_II_instruction_master_waitrequest    (nios_ii_instruction_master_waitrequest),                //                                    .waitrequest
		.nios_II_instruction_master_read           (nios_ii_instruction_master_read),                       //                                    .read
		.nios_II_instruction_master_readdata       (nios_ii_instruction_master_readdata),                   //                                    .readdata
		.memory_s1_address                         (mm_interconnect_0_memory_s1_address),                   //                           memory_s1.address
		.memory_s1_write                           (mm_interconnect_0_memory_s1_write),                     //                                    .write
		.memory_s1_readdata                        (mm_interconnect_0_memory_s1_readdata),                  //                                    .readdata
		.memory_s1_writedata                       (mm_interconnect_0_memory_s1_writedata),                 //                                    .writedata
		.memory_s1_byteenable                      (mm_interconnect_0_memory_s1_byteenable),                //                                    .byteenable
		.memory_s1_chipselect                      (mm_interconnect_0_memory_s1_chipselect),                //                                    .chipselect
		.memory_s1_clken                           (mm_interconnect_0_memory_s1_clken),                     //                                    .clken
		.nios_II_debug_mem_slave_address           (mm_interconnect_0_nios_ii_debug_mem_slave_address),     //             nios_II_debug_mem_slave.address
		.nios_II_debug_mem_slave_write             (mm_interconnect_0_nios_ii_debug_mem_slave_write),       //                                    .write
		.nios_II_debug_mem_slave_read              (mm_interconnect_0_nios_ii_debug_mem_slave_read),        //                                    .read
		.nios_II_debug_mem_slave_readdata          (mm_interconnect_0_nios_ii_debug_mem_slave_readdata),    //                                    .readdata
		.nios_II_debug_mem_slave_writedata         (mm_interconnect_0_nios_ii_debug_mem_slave_writedata),   //                                    .writedata
		.nios_II_debug_mem_slave_byteenable        (mm_interconnect_0_nios_ii_debug_mem_slave_byteenable),  //                                    .byteenable
		.nios_II_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_ii_debug_mem_slave_waitrequest), //                                    .waitrequest
		.nios_II_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_ii_debug_mem_slave_debugaccess)  //                                    .debugaccess
	);

	processor_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (nios_ii_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_ii_debug_reset_request_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
