module Component (
	dataa,
	result,
	led
);

input dataa;
output result;
output wire led;

assign result = led;
assign led = 0;

endmodule

