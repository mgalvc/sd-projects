// nios.v

// Generated using ACDS version 13.1 162 at 2018.10.05.14:27:30

`timescale 1 ps / 1 ps
module nios (
		input  wire       clk_clk,                         //                      clk.clk
		input  wire       reset_reset_n,                   //                    reset.reset_n
		input  wire [3:0] buttons_connection_export,       //       buttons_connection.export
		output wire [4:0] leds_connection_export,          //          leds_connection.export
		output wire       lcd_rs_export,                   //                   lcd_rs.export
		output wire       lcd_rw_export,                   //                   lcd_rw.export
		output wire [7:0] lcd_data_export,                 //                 lcd_data.export
		output wire       lcd_en_export,                   //                   lcd_en.export
		output wire       lcd_custom_0_conduit_end_export  // lcd_custom_0_conduit_end.export
	);

	wire  [31:0] nios2_custom_instruction_master_result;                                  // nios2_custom_instruction_master_translator:ci_slave_result -> nios2:E_ci_result
	wire   [4:0] nios2_custom_instruction_master_b;                                       // nios2:D_ci_b -> nios2_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_custom_instruction_master_c;                                       // nios2:D_ci_c -> nios2_custom_instruction_master_translator:ci_slave_c
	wire   [4:0] nios2_custom_instruction_master_a;                                       // nios2:D_ci_a -> nios2_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] nios2_custom_instruction_master_n;                                       // nios2:D_ci_n -> nios2_custom_instruction_master_translator:ci_slave_n
	wire         nios2_custom_instruction_master_writerc;                                 // nios2:D_ci_writerc -> nios2_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_dataa;                                   // nios2:E_ci_dataa -> nios2_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_custom_instruction_master_readra;                                  // nios2:D_ci_readra -> nios2_custom_instruction_master_translator:ci_slave_readra
	wire  [31:0] nios2_custom_instruction_master_datab;                                   // nios2:E_ci_datab -> nios2_custom_instruction_master_translator:ci_slave_datab
	wire         nios2_custom_instruction_master_readrb;                                  // nios2:D_ci_readrb -> nios2_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios2_custom_instruction_master_translator_comb_ci_master_result;        // nios2_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_custom_instruction_master_translator:comb_ci_master_result
	wire   [4:0] nios2_custom_instruction_master_translator_comb_ci_master_b;             // nios2_custom_instruction_master_translator:comb_ci_master_b -> nios2_custom_instruction_master_comb_xconnect:ci_slave_b
	wire   [4:0] nios2_custom_instruction_master_translator_comb_ci_master_c;             // nios2_custom_instruction_master_translator:comb_ci_master_c -> nios2_custom_instruction_master_comb_xconnect:ci_slave_c
	wire  [31:0] nios2_custom_instruction_master_translator_comb_ci_master_dataa;         // nios2_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire   [4:0] nios2_custom_instruction_master_translator_comb_ci_master_a;             // nios2_custom_instruction_master_translator:comb_ci_master_a -> nios2_custom_instruction_master_comb_xconnect:ci_slave_a
	wire         nios2_custom_instruction_master_translator_comb_ci_master_readra;        // nios2_custom_instruction_master_translator:comb_ci_master_readra -> nios2_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [7:0] nios2_custom_instruction_master_translator_comb_ci_master_n;             // nios2_custom_instruction_master_translator:comb_ci_master_n -> nios2_custom_instruction_master_comb_xconnect:ci_slave_n
	wire         nios2_custom_instruction_master_translator_comb_ci_master_writerc;       // nios2_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_translator_comb_ci_master_datab;         // nios2_custom_instruction_master_translator:comb_ci_master_datab -> nios2_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_translator_comb_ci_master_ipending;      // nios2_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire         nios2_custom_instruction_master_translator_comb_ci_master_readrb;        // nios2_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire         nios2_custom_instruction_master_translator_comb_ci_master_estatus;       // nios2_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_result;         // nios2_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_custom_instruction_master_comb_xconnect:ci_master0_result
	wire   [4:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_b;              // nios2_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire   [4:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_c;              // nios2_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire  [31:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // nios2_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire   [4:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_a;              // nios2_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire         nios2_custom_instruction_master_comb_xconnect_ci_master0_readra;         // nios2_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [7:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_n;              // nios2_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire         nios2_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // nios2_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_datab;          // nios2_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // nios2_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire         nios2_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // nios2_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire         nios2_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // nios2_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_custom_instruction_master_comb_slave_translator0_ci_master_result; // LCD_Custom_0:result -> nios2_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // nios2_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> LCD_Custom_0:dataa
	wire  [31:0] mm_interconnect_0_lcd_rw_s1_writedata;                                   // mm_interconnect_0:lcd_rw_s1_writedata -> lcd_rw:writedata
	wire   [1:0] mm_interconnect_0_lcd_rw_s1_address;                                     // mm_interconnect_0:lcd_rw_s1_address -> lcd_rw:address
	wire         mm_interconnect_0_lcd_rw_s1_chipselect;                                  // mm_interconnect_0:lcd_rw_s1_chipselect -> lcd_rw:chipselect
	wire         mm_interconnect_0_lcd_rw_s1_write;                                       // mm_interconnect_0:lcd_rw_s1_write -> lcd_rw:write_n
	wire  [31:0] mm_interconnect_0_lcd_rw_s1_readdata;                                    // lcd_rw:readdata -> mm_interconnect_0:lcd_rw_s1_readdata
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                     // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                       // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                    // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire         mm_interconnect_0_leds_s1_write;                                         // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                      // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                    // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                      // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                        // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                          // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                           // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                       // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_lcd_en_s1_writedata;                                   // mm_interconnect_0:lcd_en_s1_writedata -> lcd_en:writedata
	wire   [1:0] mm_interconnect_0_lcd_en_s1_address;                                     // mm_interconnect_0:lcd_en_s1_address -> lcd_en:address
	wire         mm_interconnect_0_lcd_en_s1_chipselect;                                  // mm_interconnect_0:lcd_en_s1_chipselect -> lcd_en:chipselect
	wire         mm_interconnect_0_lcd_en_s1_write;                                       // mm_interconnect_0:lcd_en_s1_write -> lcd_en:write_n
	wire  [31:0] mm_interconnect_0_lcd_en_s1_readdata;                                    // lcd_en:readdata -> mm_interconnect_0:lcd_en_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                                    // mm_interconnect_0:buttons_s1_address -> buttons:address
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                                   // buttons:readdata -> mm_interconnect_0:buttons_s1_readdata
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                                   // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire  [10:0] mm_interconnect_0_memory_s1_address;                                     // mm_interconnect_0:memory_s1_address -> memory:address
	wire         mm_interconnect_0_memory_s1_chipselect;                                  // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire         mm_interconnect_0_memory_s1_clken;                                       // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_memory_s1_write;                                       // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                                    // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                                  // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;                   // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;                     // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;                       // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;                         // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;                          // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;                      // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;                   // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;                    // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire         nios2_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [13:0] nios2_instruction_master_address;                                        // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                           // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                                       // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_data_master_waitrequest;                                           // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                             // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [13:0] nios2_data_master_address;                                               // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                                 // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                                  // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                              // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                                           // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire   [3:0] nios2_data_master_byteenable;                                            // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire  [31:0] mm_interconnect_0_lcd_data_s1_writedata;                                 // mm_interconnect_0:lcd_data_s1_writedata -> lcd_data:writedata
	wire   [1:0] mm_interconnect_0_lcd_data_s1_address;                                   // mm_interconnect_0:lcd_data_s1_address -> lcd_data:address
	wire         mm_interconnect_0_lcd_data_s1_chipselect;                                // mm_interconnect_0:lcd_data_s1_chipselect -> lcd_data:chipselect
	wire         mm_interconnect_0_lcd_data_s1_write;                                     // mm_interconnect_0:lcd_data_s1_write -> lcd_data:write_n
	wire  [31:0] mm_interconnect_0_lcd_data_s1_readdata;                                  // lcd_data:readdata -> mm_interconnect_0:lcd_data_s1_readdata
	wire  [31:0] mm_interconnect_0_lcd_rs_s1_writedata;                                   // mm_interconnect_0:lcd_rs_s1_writedata -> lcd_rs:writedata
	wire   [1:0] mm_interconnect_0_lcd_rs_s1_address;                                     // mm_interconnect_0:lcd_rs_s1_address -> lcd_rs:address
	wire         mm_interconnect_0_lcd_rs_s1_chipselect;                                  // mm_interconnect_0:lcd_rs_s1_chipselect -> lcd_rs:chipselect
	wire         mm_interconnect_0_lcd_rs_s1_write;                                       // mm_interconnect_0:lcd_rs_s1_write -> lcd_rs:write_n
	wire  [31:0] mm_interconnect_0_lcd_rs_s1_readdata;                                    // lcd_rs:readdata -> mm_interconnect_0:lcd_rs_s1_readdata
	wire         irq_mapper_receiver0_irq;                                                // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_d_irq_irq;                                                         // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [buttons:reset_n, irq_mapper:reset, jtag:rst_n, lcd_data:reset_n, lcd_en:reset_n, lcd_rs:reset_n, lcd_rw:reset_n, leds:reset_n, memory:reset, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, nios2:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [memory:reset_req, nios2:reset_req, rst_translator:reset_req_in]
	wire         nios2_jtag_debug_module_reset_reset;                                     // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_result                           (nios2_custom_instruction_master_result),                // custom_instruction_master.result
		.D_ci_a                                (nios2_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (nios2_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (nios2_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (nios2_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (nios2_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (nios2_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (nios2_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (nios2_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (nios2_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (),                                                      //                          .clk
		.E_ci_multi_reset                      (),                                                      //                          .reset
		.E_ci_multi_reset_req                  ()                                                       //                          .reset_req
	);

	nios_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)      //       .reset_req
	);

	nios_buttons buttons (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_buttons_s1_readdata), //                    .readdata
		.in_port  (buttons_connection_export)              // external_connection.export
	);

	nios_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_connection_export)                // external_connection.export
	);

	nios_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	nios_lcd_rs lcd_rs (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd_rs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_rs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_rs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_rs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_rs_s1_readdata),   //                    .readdata
		.out_port   (lcd_rs_export)                           // external_connection.export
	);

	nios_lcd_rs lcd_rw (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd_rw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_rw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_rw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_rw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_rw_s1_readdata),   //                    .readdata
		.out_port   (lcd_rw_export)                           // external_connection.export
	);

	nios_lcd_data lcd_data (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_lcd_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_data_s1_readdata),   //                    .readdata
		.out_port   (lcd_data_export)                           // external_connection.export
	);

	nios_lcd_rs lcd_en (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_en_s1_readdata),   //                    .readdata
		.out_port   (lcd_en_export)                           // external_connection.export
	);

	LCD lcd_custom_0 (
		.dataa  (nios2_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.result (nios2_custom_instruction_master_comb_slave_translator0_ci_master_result), //                              .result
		.LED    (lcd_custom_0_conduit_end_export)                                          //                   conduit_end.export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nios2_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nios2_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nios2_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nios2_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nios2_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nios2_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nios2_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nios2_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nios2_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (),                                                                   //               .ipending
		.ci_slave_estatus          (),                                                                   //               .estatus
		.comb_ci_master_dataa      (nios2_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nios2_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nios2_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nios2_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nios2_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nios2_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nios2_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nios2_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nios2_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nios2_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nios2_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                               //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                               //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                               //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                               //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                               //    (terminated)
		.ci_slave_multi_done       (),                                                                   //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                               //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                               //    (terminated)
		.ci_slave_multi_result     (),                                                                   //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                        //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                               //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                               //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                               //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                           //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                           //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                           //    (terminated)
		.multi_ci_master_clk       (),                                                                   //    (terminated)
		.multi_ci_master_reset     (),                                                                   //    (terminated)
		.multi_ci_master_clken     (),                                                                   //    (terminated)
		.multi_ci_master_reset_req (),                                                                   //    (terminated)
		.multi_ci_master_start     (),                                                                   //    (terminated)
		.multi_ci_master_done      (1'b0),                                                               //    (terminated)
		.multi_ci_master_dataa     (),                                                                   //    (terminated)
		.multi_ci_master_datab     (),                                                                   //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                               //    (terminated)
		.multi_ci_master_n         (),                                                                   //    (terminated)
		.multi_ci_master_readra    (),                                                                   //    (terminated)
		.multi_ci_master_readrb    (),                                                                   //    (terminated)
		.multi_ci_master_writerc   (),                                                                   //    (terminated)
		.multi_ci_master_a         (),                                                                   //    (terminated)
		.multi_ci_master_b         (),                                                                   //    (terminated)
		.multi_ci_master_c         ()                                                                    //    (terminated)
	);

	nios_nios2_custom_instruction_master_comb_xconnect nios2_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios2_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_result    (nios2_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_datab     (),                                                                        // (terminated)
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_clk       (),                                                                        // (terminated)
		.ci_master_clken     (),                                                                        // (terminated)
		.ci_master_reset_req (),                                                                        // (terminated)
		.ci_master_reset     (),                                                                        // (terminated)
		.ci_master_start     (),                                                                        // (terminated)
		.ci_master_done      (1'b0),                                                                    // (terminated)
		.ci_slave_clk        (1'b0),                                                                    // (terminated)
		.ci_slave_clken      (1'b0),                                                                    // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                    // (terminated)
		.ci_slave_reset      (1'b0),                                                                    // (terminated)
		.ci_slave_start      (1'b0),                                                                    // (terminated)
		.ci_slave_done       ()                                                                         // (terminated)
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                             (clk_clk),                                               //                           clock_clk.clk
		.nios2_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // nios2_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                 (nios2_data_master_address),                             //                   nios2_data_master.address
		.nios2_data_master_waitrequest             (nios2_data_master_waitrequest),                         //                                    .waitrequest
		.nios2_data_master_byteenable              (nios2_data_master_byteenable),                          //                                    .byteenable
		.nios2_data_master_read                    (nios2_data_master_read),                                //                                    .read
		.nios2_data_master_readdata                (nios2_data_master_readdata),                            //                                    .readdata
		.nios2_data_master_write                   (nios2_data_master_write),                               //                                    .write
		.nios2_data_master_writedata               (nios2_data_master_writedata),                           //                                    .writedata
		.nios2_data_master_debugaccess             (nios2_data_master_debugaccess),                         //                                    .debugaccess
		.nios2_instruction_master_address          (nios2_instruction_master_address),                      //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest      (nios2_instruction_master_waitrequest),                  //                                    .waitrequest
		.nios2_instruction_master_read             (nios2_instruction_master_read),                         //                                    .read
		.nios2_instruction_master_readdata         (nios2_instruction_master_readdata),                     //                                    .readdata
		.buttons_s1_address                        (mm_interconnect_0_buttons_s1_address),                  //                          buttons_s1.address
		.buttons_s1_readdata                       (mm_interconnect_0_buttons_s1_readdata),                 //                                    .readdata
		.jtag_avalon_jtag_slave_address            (mm_interconnect_0_jtag_avalon_jtag_slave_address),      //              jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write              (mm_interconnect_0_jtag_avalon_jtag_slave_write),        //                                    .write
		.jtag_avalon_jtag_slave_read               (mm_interconnect_0_jtag_avalon_jtag_slave_read),         //                                    .read
		.jtag_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),     //                                    .readdata
		.jtag_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),    //                                    .writedata
		.jtag_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),  //                                    .waitrequest
		.jtag_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),   //                                    .chipselect
		.lcd_data_s1_address                       (mm_interconnect_0_lcd_data_s1_address),                 //                         lcd_data_s1.address
		.lcd_data_s1_write                         (mm_interconnect_0_lcd_data_s1_write),                   //                                    .write
		.lcd_data_s1_readdata                      (mm_interconnect_0_lcd_data_s1_readdata),                //                                    .readdata
		.lcd_data_s1_writedata                     (mm_interconnect_0_lcd_data_s1_writedata),               //                                    .writedata
		.lcd_data_s1_chipselect                    (mm_interconnect_0_lcd_data_s1_chipselect),              //                                    .chipselect
		.lcd_en_s1_address                         (mm_interconnect_0_lcd_en_s1_address),                   //                           lcd_en_s1.address
		.lcd_en_s1_write                           (mm_interconnect_0_lcd_en_s1_write),                     //                                    .write
		.lcd_en_s1_readdata                        (mm_interconnect_0_lcd_en_s1_readdata),                  //                                    .readdata
		.lcd_en_s1_writedata                       (mm_interconnect_0_lcd_en_s1_writedata),                 //                                    .writedata
		.lcd_en_s1_chipselect                      (mm_interconnect_0_lcd_en_s1_chipselect),                //                                    .chipselect
		.lcd_rs_s1_address                         (mm_interconnect_0_lcd_rs_s1_address),                   //                           lcd_rs_s1.address
		.lcd_rs_s1_write                           (mm_interconnect_0_lcd_rs_s1_write),                     //                                    .write
		.lcd_rs_s1_readdata                        (mm_interconnect_0_lcd_rs_s1_readdata),                  //                                    .readdata
		.lcd_rs_s1_writedata                       (mm_interconnect_0_lcd_rs_s1_writedata),                 //                                    .writedata
		.lcd_rs_s1_chipselect                      (mm_interconnect_0_lcd_rs_s1_chipselect),                //                                    .chipselect
		.lcd_rw_s1_address                         (mm_interconnect_0_lcd_rw_s1_address),                   //                           lcd_rw_s1.address
		.lcd_rw_s1_write                           (mm_interconnect_0_lcd_rw_s1_write),                     //                                    .write
		.lcd_rw_s1_readdata                        (mm_interconnect_0_lcd_rw_s1_readdata),                  //                                    .readdata
		.lcd_rw_s1_writedata                       (mm_interconnect_0_lcd_rw_s1_writedata),                 //                                    .writedata
		.lcd_rw_s1_chipselect                      (mm_interconnect_0_lcd_rw_s1_chipselect),                //                                    .chipselect
		.leds_s1_address                           (mm_interconnect_0_leds_s1_address),                     //                             leds_s1.address
		.leds_s1_write                             (mm_interconnect_0_leds_s1_write),                       //                                    .write
		.leds_s1_readdata                          (mm_interconnect_0_leds_s1_readdata),                    //                                    .readdata
		.leds_s1_writedata                         (mm_interconnect_0_leds_s1_writedata),                   //                                    .writedata
		.leds_s1_chipselect                        (mm_interconnect_0_leds_s1_chipselect),                  //                                    .chipselect
		.memory_s1_address                         (mm_interconnect_0_memory_s1_address),                   //                           memory_s1.address
		.memory_s1_write                           (mm_interconnect_0_memory_s1_write),                     //                                    .write
		.memory_s1_readdata                        (mm_interconnect_0_memory_s1_readdata),                  //                                    .readdata
		.memory_s1_writedata                       (mm_interconnect_0_memory_s1_writedata),                 //                                    .writedata
		.memory_s1_byteenable                      (mm_interconnect_0_memory_s1_byteenable),                //                                    .byteenable
		.memory_s1_chipselect                      (mm_interconnect_0_memory_s1_chipselect),                //                                    .chipselect
		.memory_s1_clken                           (mm_interconnect_0_memory_s1_clken),                     //                                    .clken
		.nios2_jtag_debug_module_address           (mm_interconnect_0_nios2_jtag_debug_module_address),     //             nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write             (mm_interconnect_0_nios2_jtag_debug_module_write),       //                                    .write
		.nios2_jtag_debug_module_read              (mm_interconnect_0_nios2_jtag_debug_module_read),        //                                    .read
		.nios2_jtag_debug_module_readdata          (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                                    .readdata
		.nios2_jtag_debug_module_writedata         (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                                    .writedata
		.nios2_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                                    .byteenable
		.nios2_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                                    .waitrequest
		.nios2_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_jtag_debug_module_debugaccess)  //                                    .debugaccess
	);

	nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
